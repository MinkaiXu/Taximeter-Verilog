`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:46:16 04/16/2017 
// Design Name: 
// Module Name:    calculate_distance_sub 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module calculate_distance_sub(
	input clk,
	input park,
	input restart,
	inout reg[15:0]distance
    );

	
endmodule
